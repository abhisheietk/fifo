module dpram (
    clK, 
    a_port_WR,
    a_port_ADDR,
    a_port_data_IN,
    a_port_data_OUT,
    b_port_WR,
    b_port_ADDR,
    b_port_data_IN,
    b_port_data_OUT
);