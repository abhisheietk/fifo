module dpram (
    clK, 
    fifo_IN,
    fifo_OUT
    );

    parameter DATA = 16;
    parameter ADDR = 5;